module manipular_vetores( 
    input [31:0] entrada,
    output [31:0] saida );

    // insira seu código aqui

endmodule